module eth_sdram_dac(
    input                  sys_clk     ,  //FPGA外部时钟，50MHz
    input                  sys_rst_n   ,  //系统复位，低电平有效
    input                  touch_key   ,  //触摸按键输入，用于切换rd_en状态
    //以太网接口                          
    input                  eth_rxc     ,  //RGMII接收数据时钟
    input                  eth_rx_ctl  ,  //RGMII输入数据有效信号
    input       [3:0]      eth_rxd     ,  //RGMII输入数据
    output                 eth_txc     ,  //RGMII发送数据时钟    
    output                 eth_tx_ctl  ,  //RGMII输出数据有效信号
    output      [3:0]      eth_txd     ,  //RGMII输出数据          
    output                 eth_rst_n   ,  //以太网芯片复位信号，低电平有效   
    //SDRAM 
    output                 sdram_clk   ,  //SDRAM 时钟
    output                 sdram_cke   ,  //SDRAM 时钟有效
    output                 sdram_cs_n  ,  //SDRAM 片选
    output                 sdram_ras_n ,  //SDRAM 行有效
    output                 sdram_cas_n ,  //SDRAM 列有效
    output                 sdram_we_n  ,  //SDRAM 写有效
    output      [1:0]      sdram_ba    ,  //SDRAM Bank地址
    output      [1:0]      sdram_dqm   ,  //SDRAM 数据掩码
    output      [12:0]     sdram_addr  ,  //SDRAM 地址
    inout       [7:0]      sdram_data  ,  //SDRAM 数据                                          
    output                     dac_clk ,  
   
	 //DAC接口 - 10位DAC
	 output    [9:0]        dac_data_final
    );
                                                       
//wire define    
wire         rst_n                     ;  //复位信号
wire         clk_100m                  ;
wire         clk_100m_shift            ;
wire         clk_50m                   ;  //50mhz时钟
wire         clk_1m                   ;  //1mhz时钟,提供给dac驱动时钟
wire         locked                    ;  //时钟锁定信号  

wire         gmii_rx_clk               ;  //以太网125M时钟                                         
wire         rdata_req                 ;  //SDRAM控制器模块读使能
wire  [7:0] rd_data                   ;  //SDRAM控制器模块读数据
wire         sdram_init_done           ;  //SDRAM初始化完成sdram_init_done
wire  [23:0] sdram_max_addr            ;  //存入SDRAM的最大读写地址，修正为24位 
wire  [31:0] rec_data                  ;  //以太网接收的数据
wire        dac_data_req               ;
wire  [7:0] dac_data_to_controller     ;
wire        dac_data_valid             ;
wire        rec_en                     ; 
wire [7:0] sdram_rd_data              ;
wire  [7:0] dac_data                    ;
wire        rd_en_ctrl                 ;  //按键控制的读使能信号
//*****************************************************
//**                    main code
//*****************************************************

assign rst_n = sys_rst_n & locked;
//系统初始化完成：SDRAM初始化完成
//修正地址计算：8MB = 8*1024*1024 = 8388608字节
//由于突发长度为512，实际可用地址应该为 8388608 + 512 = 8389120 
//但考虑到24位地址限制，设置为8388608 + 512 = 8389120，确保完整的8MB数据可以存储
//这里根据实际DAC输出情况尝试除以4 得到2097152
assign sdram_max_addr = 24'd2097152; //8MB数据 + 突发长度补偿

//锁相环
pll_clk u_pll_clk(
    .areset             (~sys_rst_n    ),
    .inclk0             (sys_clk       ),
            
    .c0                 (clk_100m      ),
    .c1                 (clk_100m_shift),
    .c2                 (clk_50m       ),
    .c3                 (clk_1m)        ,
    .locked             (locked        )
    );
    
//以太网顶层
eth_top u_eth_top(
    .sys_rst_n          (rst_n) ,           //系统复位信号，低电平有效 
    .eth_rxc            (eth_rxc)   ,       //RGMII接收数据时钟
    .eth_rx_ctl         (eth_rx_ctl),       //RGMII输入数据有效信号
    .eth_rxd            (eth_rxd)   ,       //RGMII输入数据
    .eth_txc            (eth_txc)   ,       //RGMII发送数据时钟    
    .eth_tx_ctl         (eth_tx_ctl),       //RGMII输出数据有效信号
    .eth_txd            (eth_txd)   ,       //RGMII输出数据          
    .eth_rst_n          (eth_rst_n) ,       //以太网芯片复位信号，低电平有效 

    .rec_en             (rec_en),           //以太网32位数据接收完成
    .rec_data           (rec_data),         //以太网32位数据
    .gmii_rx_clk        (gmii_rx_clk)       //以太网125M时钟
    ); 

//触摸按键模块，用于控制SDRAM读使能
//复位时rd_en_ctrl默认为低电平，禁用SDRAM读操作
//按键按下时切换rd_en_ctrl状态
touch u_touch(
    .clk_50m            (clk_50m),          //50MHz时钟
    .rst_n              (rst_n),            //复位信号
    .touch_key          (touch_key),        //触摸按键输入
    .touch_cnt          (rd_en_ctrl)        //输出读使能控制信号
    );
    
udp_32_to_8bit u_udp_32_to_8bit(    
    .clk        (gmii_rx_clk)   ,
    .rst_n      (rst_n )      ,
    .rec_en     (rec_en)     ,   
    .rec_data   (rec_data) ,                  
    .dac_data   (dac_data_to_controller) ,                    
    .data_valid (dac_data_valid)    
);
    
//SDRAM 控制器顶层模块,封装成FIFO接口
//SDRAM 控制器地址组成: {bank_addr[1:0],row_addr[12:0],col_addr[8:0]}
sdram_top u_sdram_top(
    .ref_clk            (clk_100m),         //sdram 控制器参考时钟
    .out_clk            (clk_100m_shift),   //用于输出的相位偏移时钟
    .rst_n              (rst_n),            //系统复位
                                            
    //用户写端口                              
    .wr_clk             (gmii_rx_clk),      //写端口FIFO: 写时钟
    .wr_en              (dac_data_valid),                          //写端口FIFO: 写使能
    .wr_data            (dac_data_to_controller),         //写端口FIFO: 写数据
    .wr_min_addr        (24'd0),            //写SDRAM的起始地址
    .wr_max_addr        (sdram_max_addr),   //写SDRAM的结束地址
    .wr_len             (10'd512),          //写SDRAM时的数据突发长度
    .wr_load            (~rst_n),           //写端口复位: 复位写地址,清空写FIFO
                                            
    //用户读端口                              
    .rd_clk             (clk_1m),          //读端口FIFO: 读时钟
    .rd_en              (rd_en_ctrl),      //读端口FIFO: 读使能，由按键控制，读FIFO到DAC
    .rd_data            (sdram_rd_data),    //读端口FIFO: 读数据
    .rd_min_addr        (24'd0),            //读SDRAM的起始地址
    .rd_max_addr        (sdram_max_addr),   //读SDRAM的结束地址
    .rd_len             (10'd512),          //从SDRAM中读数据时的突发长度
    .rd_load            (~rst_n),           //读端口复位: 复位读地址,清空读FIFO
                                                
    //用户控制端口                                
    .sdram_read_valid   (1'b1),             //SDRAM 读使能  SDRAM进读FIFO
    .sdram_pingpang_en  (1'b0),             //SDRAM 乒乓操作使能
    .sdram_init_done    (sdram_init_done),  //SDRAM 初始化完成标志
                                            
    //SDRAM 芯片接口                                
    .sdram_clk          (sdram_clk),        //SDRAM 芯片时钟
    .sdram_cke          (sdram_cke),        //SDRAM 时钟有效
    .sdram_cs_n         (sdram_cs_n),       //SDRAM 片选
    .sdram_ras_n        (sdram_ras_n),      //SDRAM 行有效
    .sdram_cas_n        (sdram_cas_n),      //SDRAM 列有效
    .sdram_we_n         (sdram_we_n),       //SDRAM 写有效
    .sdram_ba           (sdram_ba),         //SDRAM Bank地址
    .sdram_addr         (sdram_addr),       //SDRAM 行/列地址
    .sdram_data         (sdram_data),       //SDRAM 数据
    .sdram_dqm          (sdram_dqm)         //SDRAM 数据掩码
    );



assign dac_clk = clk_50m;


//10BIT-DAC使用： 直接使用8位数据，末端2位补0
assign dac_data_final = {sdram_rd_data,2'b0};    //8位+2位0

endmodule 